library verilog;
use verilog.vl_types.all;
entity compare_8bit_vlg_vec_tst is
end compare_8bit_vlg_vec_tst;
