library verilog;
use verilog.vl_types.all;
entity upcounter_vlg_vec_tst is
end upcounter_vlg_vec_tst;
