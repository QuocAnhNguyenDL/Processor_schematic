library verilog;
use verilog.vl_types.all;
entity sel8to1_8bit_vlg_vec_tst is
end sel8to1_8bit_vlg_vec_tst;
