library verilog;
use verilog.vl_types.all;
entity compare_8bit_vlg_check_tst is
    port(
        less            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end compare_8bit_vlg_check_tst;
