library verilog;
use verilog.vl_types.all;
entity downcounter_vlg_vec_tst is
end downcounter_vlg_vec_tst;
