library verilog;
use verilog.vl_types.all;
entity sel4to1_8bit_vlg_vec_tst is
end sel4to1_8bit_vlg_vec_tst;
