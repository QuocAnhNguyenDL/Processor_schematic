library verilog;
use verilog.vl_types.all;
entity Dmem_vlg_vec_tst is
end Dmem_vlg_vec_tst;
