library verilog;
use verilog.vl_types.all;
entity sel8to1_8bit_vlg_check_tst is
    port(
        R               : in     vl_logic_vector(7 downto 0);
        sampler_rx      : in     vl_logic
    );
end sel8to1_8bit_vlg_check_tst;
